module mojo_top(
    // 50MHz clock input
    input clk,
    // Input from reset button (active low)
    input rst_n,
    // cclk input from AVR, high when AVR is ready
    input cclk,
    // Outputs to the 8 onboard LEDs
    output[7:0]led,
    // AVR SPI connections
    output spi_miso,
    input spi_ss,
    input spi_mosi,
    input spi_sck,
    // AVR ADC channel select
    output [3:0] spi_channel,
    // Serial connections
    input avr_tx, // AVR Tx => FPGA Rx
    output avr_rx, // AVR Rx => FPGA Tx
    input avr_rx_busy // AVR Rx buffer full
    );

wire rst = ~rst_n; // make reset active high

// these signals should be high-z when not used
assign spi_miso = 1'bz;
assign avr_rx = 1'bz;
assign spi_channel = 4'bzzzz;

microblaze_mcs mcs_0 (
	.Clk(clk), // input Clk
	.Reset(rst), // input Reset
	.FIT1_Interrupt(), // output FIT1_Interrupt
	.FIT1_Toggle(), // output FIT1_Toggle
	.GPO1(led), // output [7 : 0] GP01
	.INTC_IRQ() // output INTC_IRQ
);

endmodule